
module Flash_loader (
	noe_in);	

	input		noe_in;
endmodule
