module omdazz_cyclon_iv_devoard_top
(
    
);

endmodule
