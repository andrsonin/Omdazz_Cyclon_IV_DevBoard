// altclkctrl_inst.v

// Generated using ACDS version 22.1 915

`timescale 1 ps / 1 ps
module altclkctrl_inst (
		input  wire  inclk,  //  altclkctrl_input.inclk
		input  wire  ena,    //                  .ena
		output wire  outclk  // altclkctrl_output.outclk
	);

	Flash_loader_serial_flash_loader_0_altclkctrl_inst_altclkctrl_inst altclkctrl_inst (
		.inclk  (inclk),  //  altclkctrl_input.inclk
		.ena    (ena),    //                  .ena
		.outclk (outclk)  // altclkctrl_output.outclk
	);

endmodule
